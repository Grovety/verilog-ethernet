module phytest (
);

endmodule
