module phytest
(
);
endmodule
